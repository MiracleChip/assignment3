`timescale 1ns/1ps
`define NUM_FLOORS 10                    // Number of floors
`define FLOOR_BITS $clog2(`NUM_FLOORS)    // Bits to represent the number of floors
